module line_state_detector_tb ();
endmodule